module this_module (
    input i_1,
    input i_2,
    output o_1,
);

    assign o_1 = i_1 | i_2;

endmodule